module cla_64bit( a, b, cin, sum, cout);

	input [63:0] a, b;
	input cin;
	output [63:0] sum;
	output cout;
	//write your design below

	
endmodule



